//-------------------------------------------------------------------------------------------------
module saa1099
//-------------------------------------------------------------------------------------------------
(
	input  wire      clk_sys,
	input  wire      ce,      // 8 MHz
	input  wire      rst_n,
	input  wire      cs_n,
	input  wire      a0,      // 0=data, 1=address
	input  wire      wr_n,
	input  wire[7:0] din,
	output wire[7:0] out_r,
	output wire[7:0] out_l
);
//-------------------------------------------------------------------------------------------------

assign out_r = 8'd0;
assign out_l = 8'd0;

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
