//-------------------------------------------------------------------------------------------------
module specdrum
//-------------------------------------------------------------------------------------------------
(
	input  wire      clock,
	input  wire      ce,
	input  wire      iorq,
	input  wire      wr,
	input  wire[7:0] d,
	output reg [7:0] q,
	input  wire[7:4] a
);
//-------------------------------------------------------------------------------------------------

always @(posedge clock) if(ce) if(!iorq && !wr && a == 4'b1101) q <= d;

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
