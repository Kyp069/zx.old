//-------------------------------------------------------------------------------------------------
module clock
//-------------------------------------------------------------------------------------------------
(
	input  wire       i,
	input  wire       model,
	output wire       clock,
	output wire       power,

	output reg        ne14M,

	output reg        pe7M0,
	output reg        ne7M0,

	output reg        pe3M5,
	output reg        ne3M5
);
//-------------------------------------------------------------------------------------------------

wire ci;
IBUFG IBufg(.I(i), .O(ci));

//-------------------------------------------------------------------------------------------------

wire b0, c0, l0, o0;

DCM_SP #
(
	.CLKIN_PERIOD          (20.000),
	.CLKDV_DIVIDE          ( 2.000),
	.CLKFX_DIVIDE          (25    ),
	.CLKFX_MULTIPLY        (28    )
)
Dcm0
(
	.RST                   (1'b0),
	.DSSEN                 (1'b0),
	.PSCLK                 (1'b0),
	.PSEN                  (1'b0),
	.PSINCDEC              (1'b0),
	.CLKIN                 (ci),
	.CLKFB                 (b0),
	.CLK0                  (c0),
	.CLK90                 (),
	.CLK180                (),
	.CLK270                (),
	.CLK2X                 (),
	.CLK2X180              (),
	.CLKFX                 (o0), // 56.000 MHz output
	.CLKFX180              (),
	.CLKDV                 (),
	.PSDONE                (),
	.STATUS                (),
	.LOCKED                (l0)
);

BUFG Bufg0(.I(c0), .O(b0));

//-------------------------------------------------------------------------------------------------

wire b1, c1, l1, o1;

DCM_SP #
(
	.CLKIN_PERIOD          (20.000),
	.CLKDV_DIVIDE          ( 2.000),
	.CLKFX_DIVIDE          (22    ),
	.CLKFX_MULTIPLY        (25    )
)
Dcm1
(
	.RST                   (1'b0),
	.DSSEN                 (1'b0),
	.PSCLK                 (1'b0),
	.PSEN                  (1'b0),
	.PSINCDEC              (1'b0),
	.CLKIN                 (ci),
	.CLKFB                 (b1),
	.CLK0                  (c1),
	.CLK90                 (),
	.CLK180                (),
	.CLK270                (),
	.CLK2X                 (),
	.CLK2X180              (),
	.CLKFX                 (o1), // 56.7504 MHz output
	.CLKFX180              (),
	.CLKDV                 (),
	.PSDONE                (),
	.STATUS                (),
	.LOCKED                (l1)
);

BUFG Bufg1(.I(c1), .O(b1));

//-------------------------------------------------------------------------------------------------

BUFGMUX_1 BufgMux(.I0(o0), .I1(o1), .O(clock), .S(model));

//-------------------------------------------------------------------------------------------------

reg[3:0] ce = 4'd1;
always @(negedge clock) if(power) begin
	ce <= ce+1'd1;
	ne14M <= ~ce[0] & ~ce[1];
	pe7M0 <= ~ce[0] & ~ce[1] &  ce[2];
	ne7M0 <= ~ce[0] & ~ce[1] & ~ce[2];
	pe3M5 <= ~ce[0] & ~ce[1] & ~ce[2] &  ce[3];
	ne3M5 <= ~ce[0] & ~ce[1] & ~ce[2] & ~ce[3];
end

//-------------------------------------------------------------------------------------------------

assign power = l0 & l1;

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
